module master(
    input  wire        ACLK,
    input  wire        ARESETn,

    // Write Address
    output reg  [31:0] M_AXI_AWADDR,
    output reg         M_AXI_AWVALID,
    input  wire        M_AXI_AWREADY,
    output reg  [2:0]  M_AXI_AWPROT,

    output reg  [3:0]  M_AXI_AWID,
    output reg  [7:0]  M_AXI_AWLEN,
    output reg  [2:0]  M_AXI_AWSIZE,
    output reg  [1:0]  M_AXI_AWBURST,

    output reg  [3:0]  M_AXI_AWCACHE,
    output reg         M_AXI_AWLOCK,
    output reg  [3:0]  M_AXI_AWQOS,
    output reg  [3:0]  M_AXI_AWREGION,

    // Write Data
    output reg  [31:0] M_AXI_WDATA,
    output reg  [3:0]  M_AXI_WSTRB,
    output reg         M_AXI_WVALID,
    input  wire        M_AXI_WREADY,

    output reg         M_AXI_WLAST,

    // Write Response
    input  wire [1:0]  M_AXI_BRESP,
    input  wire        M_AXI_BVALID,
    output reg         M_AXI_BREADY,

    input  wire [3:0]  M_AXI_BID,

    // Read Address
    output reg  [31:0] M_AXI_ARADDR,
    output reg         M_AXI_ARVALID,
    input  wire        M_AXI_ARREADY,
    output reg  [2:0]  M_AXI_ARPROT,

    output reg  [3:0]  M_AXI_ARID,
    output reg  [7:0]  M_AXI_ARLEN,
    output reg  [2:0]  M_AXI_ARSIZE,
    output reg  [1:0]  M_AXI_ARBURST,

    output reg  [3:0]  M_AXI_ARCACHE,
    output reg         M_AXI_ARLOCK,
    output reg  [3:0]  M_AXI_ARQOS,
    output reg  [3:0]  M_AXI_ARREGION,

    // Read Data
    input  wire [31:0] M_AXI_RDATA,
    input  wire [1:0]  M_AXI_RRESP,
    input  wire        M_AXI_RVALID,
    output reg         M_AXI_RREADY,

    input  wire [3:0]  M_AXI_RID,
    input  wire        M_AXI_RLAST
);

parameter RESET_WAIT = 0, RUN = 1, DONE = 2;
reg [1:0] state;

// burst
localparam BURST_LEN = 4;       // beats
reg [7:0] w_beat_cnt;           // beat count of current burst

// outstanding
localparam TOTAL_BURSTS = 8;
localparam MAX_WR_OUTSTANDING = 2;
reg [2:0] wr_outstanding;       // not yet response number
reg [7:0] bursts_left;          // how many burst left (TOTAL_BURSTS)
reg sending_w;                  // whether sending w burst now

wire can_issue;
assign can_issue = 
    (bursts_left > 0) && 
    (wr_outstanding < MAX_WR_OUTSTANDING) && 
    !M_AXI_AWVALID && 
    !sending_w;

always @(posedge ACLK) begin
    if (!ARESETn) begin
        state <= RESET_WAIT;

        // AW
        M_AXI_AWVALID <= 0;
        M_AXI_AWPROT <= 0;
        M_AXI_AWID <= 0;
        M_AXI_AWLEN <= 0;
        M_AXI_AWSIZE <= 3'b010;
        M_AXI_AWBURST <= 2'b01;
        M_AXI_AWCACHE <= 4'b0011;
        M_AXI_AWLOCK <= 0;
        M_AXI_AWQOS <= 0;
        M_AXI_AWREGION <= 0;

        // W
        M_AXI_WVALID  <= 0;
        M_AXI_WLAST <= 0;

        // B
        M_AXI_BREADY  <= 1;         // always ready !!!

        // outstanding
        bursts_left <= TOTAL_BURSTS;
        sending_w <= 0;

        // AR
        M_AXI_ARVALID <= 0;
        M_AXI_ARPROT <= 0;
        M_AXI_ARID    <= 0;
        M_AXI_ARLEN   <= 0;
        M_AXI_ARSIZE  <= 3'b010;
        M_AXI_ARBURST <= 2'b01;
        M_AXI_ARCACHE <= 4'b0011;
        M_AXI_ARLOCK <= 0;
        M_AXI_ARQOS <= 0;
        M_AXI_ARREGION <= 0;

        // R
        M_AXI_RREADY  <= 0;
    end else begin
        case (state)
            RESET_WAIT: begin
                state <= RUN;
            end
            RUN: begin
                // Issue new AW
                if (can_issue) begin
                    M_AXI_AWADDR  <= 32'h0000_0000 + (TOTAL_BURSTS - bursts_left) * 16;
                    M_AXI_AWLEN   <= BURST_LEN - 1;
                    M_AXI_AWSIZE  <= 3'b010;
                    M_AXI_AWBURST <= 2'b01;
                    M_AXI_AWVALID <= 1;

                    // start W burst
                    sending_w <= 1;
                    w_beat_cnt <= 0;

                    M_AXI_WDATA <= 32'h1000_0000 + (TOTAL_BURSTS - bursts_left) * 16;
                    M_AXI_WSTRB <= 4'b1111;
                    M_AXI_WVALID<= 1;
                    M_AXI_WLAST <= 0;

                    bursts_left <= bursts_left - 1;
                end 

                // AW handshake
                if (M_AXI_AWVALID && M_AXI_AWREADY) begin
                    M_AXI_AWVALID <= 0;
                end

                // W channel
                if (sending_w && M_AXI_WVALID && M_AXI_WREADY) begin
                    w_beat_cnt <= w_beat_cnt + 1;
                    M_AXI_WDATA <= M_AXI_WDATA + 1;

                    if (w_beat_cnt == BURST_LEN - 2) begin
                        M_AXI_WLAST <= 1;
                    end
                    else if (w_beat_cnt == BURST_LEN - 1) begin
                        M_AXI_WVALID <= 0;
                        M_AXI_WLAST  <= 0;
                        sending_w    <= 0;
                    end
                end

                if ((bursts_left == 0) && (wr_outstanding == 0) && !sending_w && !M_AXI_AWVALID) begin
                    state <= DONE;
                end 
            end
            DONE: begin
                state <= DONE;
            end
        endcase
    end
end

// Independent B channel
always @(posedge ACLK) begin
    if (!ARESETn) begin
        wr_outstanding <= 0;
    end else begin
        case ({M_AXI_AWVALID && M_AXI_AWREADY,
               M_AXI_BVALID  && M_AXI_BREADY})
            2'b10: wr_outstanding <= wr_outstanding + 1;
            2'b01: wr_outstanding <= wr_outstanding - 1;
            2'b11: wr_outstanding <= wr_outstanding; // same cycle issue + complete
            default: wr_outstanding <= wr_outstanding;
        endcase
    end
end

endmodule
